library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY VGA IS
PORT(
	CLOCK_50: 				IN STD_LOGIC; --SYSTEM CLOCK
	VGA_HS, VGA_VS: 		OUT STD_LOGIC; -- HORIZONTAL AND VERTICAL SYNCRONIZATION
	VGA_R, VGA_G, VGA_B: OUT STD_LOGIC_VECTOR(7 downto 0); -- COLORS
	VGA_CLOCK:				OUT STD_LOGIC;	-- VGA CLOCK OUT
	
	KEYB_CLOCK:				IN STD_LOGIC;
	KEYDATA:					IN STD_LOGIC
);
END VGA;

ARCHITECTURE MAIN OF VGA IS


	SIGNAL VGACLK, RESET:	STD_LOGIC := '0';
	
	------------------------------

	-- PLL
	COMPONENT PLL IS
	PORT(
		CLK_IN_CLK:		IN 	STD_LOGIC := 'X'; --CLK
		RESET_RESET:	IN 	STD_LOGIC := 'X'; --RESET
		CLK_OUT_CLK:	OUT 	STD_LOGIC
	);
	END COMPONENT PLL;
	
	------------------------------
	
	-- SYN
	COMPONENT SYNC IS
	PORT(
		CLK:				IN 	STD_LOGIC; --PLL
		HSYNC, VSYNC:	OUT 	STD_LOGIC;
		R, G, B:			OUT 	STD_LOGIC_VECTOR(7 downto 0);
		CLK_KEYBOARD:	IN STD_LOGIC;
		DATA_KEY:		IN STD_LOGIC;
		CLK_50:			IN STD_LOGIC
	);
	END COMPONENT SYNC;
	
BEGIN
	C1: SYNC PORT MAP(VGACLK, VGA_HS, VGA_VS, VGA_R, VGA_G, VGA_B, KEYB_CLOCK, KEYDATA, CLOCK_50);
	C2: PLL PORT MAP(CLOCK_50, RESET, VGACLK);
	VGA_CLOCK <= VGACLK;
END MAIN;