library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY VGA IS
PORT(
	CLOCK_50: 				IN STD_LOGIC; --SYSTEM CLOCK
	VGA_HS, VGA_VS: 		OUT STD_LOGIC; -- HORIZONTAL AND VERTICAL SYNCRONIZATION
	VGA_R, VGA_G, VGA_B: OUT STD_LOGIC_VECTOR(7 downto 0); -- COLORS
	VGA_CLOCK:				OUT STD_LOGIC;	-- VGA CLOCK OUT
	
	PS2_CLK:	 IN STD_LOGIC;
	PS2_DATA: IN STD_LOGIC
);
END VGA;

ARCHITECTURE MAIN OF VGA IS


	SIGNAL VGACLK, RESET:	STD_LOGIC := '0';

	-- PLL
	COMPONENT PLL IS
	PORT(
		CLK_IN_CLK:		IN 	STD_LOGIC := 'X'; --CLK
		RESET_RESET:	IN 	STD_LOGIC := 'X'; --RESET
		CLK_OUT_CLK:	OUT 	STD_LOGIC
	);
	END COMPONENT PLL;
	
	-- SYNC
	COMPONENT SYNC IS
	PORT(
		CLK:				IN 	STD_LOGIC; --PLL
		HSYNC, VSYNC:	OUT 	STD_LOGIC;
		R, G, B:			OUT 	STD_LOGIC_VECTOR(7 downto 0)
	);
	END COMPONENT SYNC;
	
	-- KEYBOARD COMPONENT 
	COMPONENT keyboard IS
		PORT(
			clk_keyboard: IN 	STD_LOGIC; -- Pin used to emulate the clk_keyboard cycles
			data: 			IN 	STD_LOGIC	 -- Pin used for data input 
		);
	END COMPONENT keyboard;
	
	
	
BEGIN
	C1: SYNC PORT MAP(VGACLK, VGA_HS, VGA_VS, VGA_R, VGA_G, VGA_B);
	C2: PLL PORT MAP(CLOCK_50, RESET, VGACLK);
	C3:	keyboard PORT MAP(PS2_CLK, PS2_DATA);
	VGA_CLOCK <= VGACLK;
END MAIN;